library IEEE;
use IEEE.std_logic_1164.all;

entity decod_3_8 is
    port (
        sel    : in std_logic_vector (2 downto 0);
        hab    : in std_logic;
        salida : out std_logic_vector (7 downto 0));
end decod_3_8;

architecture solucion of decod_3_8 is
begin
-- Escribe aquí tu solución.
end solucion;

