library IEEE;
use IEEE.std_logic_1164.all;

entity decod_2_4 is
    port (
        sel    : in std_logic_vector (1 downto 0);
        hab    : in std_logic;
        salida : out std_logic_vector (3 downto 0));
end decod_2_4;

architecture solucion of decod_2_4 is
begin
-- Escribe aquí tu solución.
end solucion;

