library IEEE;
use IEEE.std_logic_1164.all;
use work.tp8.all;

entity cod_8_3 is
    port (
        entrada : in std_logic_vector (7 downto 0);
        valido  : out std_logic;
        salida  : out std_logic_vector (2 downto 0));
end cod_8_3;

architecture solucion of cod_8_3 is
begin
-- Escribe aquí tu solución.
end solucion;

